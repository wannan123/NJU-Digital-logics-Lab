module segs (
    input reg [7:0] ledr,
    output [7:0] seg0,
    output [7:0] seg1);
    
always @ (ledr[3:0]) begin
	case(ledr[3:0])
		4'b0000: seg0 = 8'b00000010;
		4'b0001: seg0 = 8'b10011111;
		4'b0010: seg0 = 8'b00100101;
		4'b0011: seg0 = 8'b00001101;
		4'b0100: seg0 = 8'b10011001;
		4'b0101: seg0 = 8'b01001001;
		4'b0110: seg0 = 8'b01000001;
		4'b0111: seg0 = 8'b00011111;
		4'b1000: seg0 = 8'b00000001;
		4'b1001: seg0 = 8'b00011001;
		4'b1010: seg0 = 8'b00010001;
		4'b1011: seg0 = 8'b11000001;
		4'b1100: seg0 = 8'b01100011;
		4'b1101: seg0 = 8'b10000101;
		4'b1110: seg0 = 8'b01100001;
		4'b1111: seg0 = 8'b01110001;
		default seg0 = 8'b00000010;
	endcase
end

always @ (ledr[7:4]) begin
	case(ledr[7:4])
		4'b0000: seg1 = 8'b00000010;
		4'b0001: seg1 = 8'b10011111;
		4'b0010: seg1 = 8'b00100101;
		4'b0011: seg1 = 8'b00001101;
		4'b0100: seg1 = 8'b10011001;
		4'b0101: seg1 = 8'b01001001;
		4'b0110: seg1 = 8'b01000001;
		4'b0111: seg1 = 8'b00011111;
		4'b1000: seg1 = 8'b00000001;
		4'b1001: seg1 = 8'b00011001;
		4'b1010: seg1 = 8'b00010001;
		4'b1011: seg1 = 8'b11000001;
		4'b1100: seg1 = 8'b01100011;
		4'b1101: seg1 = 8'b10000101;
		4'b1110: seg1 = 8'b01100001;
		4'b1111: seg1 = 8'b01110001;
		default seg1 = 8'b00000010;
	endcase
end
endmodule
